module Counter
(
	input clk, countStartTrigger,
	output countValue, Frequency

);

endmodule